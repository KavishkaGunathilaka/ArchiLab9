library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.numeric_std.all ;

entity ent is
  port (
    clock
  ) ;
end ent ; 

architecture arch of ent is

begin

end architecture ;